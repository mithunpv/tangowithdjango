b0VIM 7.3      ��W�k ��  mithun                                  angarr.local                            ~mithun/tangowithdjango/rango/views.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                                   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad  1   }     �       �  �  W  0    �  �  �  �  �  �  �  �  l  D  /    �  �  �  �  h  =  )  �  �  �  �  8  7  6  5  !  �  �  �  �  �  �  �  �  �  `  4  �
  �
  �
  �
  �
  l
  k
  j
  i
  T
  P
  '
  &
  %
  
  �	  �	  �	  �	  �	  �	  �	  t	  h	  @	  ,	  	  �  �  �  �  p  Q              �  �  �  �  �  �  �  �  x  l  P  3    �  �  �  �  �  |  p  K  '    
  �  �  �  �  �  e  T  4    �    Z  I  G  	  �  �  �  �  �  �  �  �  `  J  2    �  �  �  �  �  }  |                                                   			message=cd['message'] 			name=cd['name'] 				toemail=['noreply@example.com'] 			else: 				toemail=[cd['email'],]         		if cd['email']: 			fromemail=settings.EMAIL_HOST_USER; 			cd=form.cleaned_data 		if form.is_valid(): 		form=ContactForm(request.POST) 	if request.method=='POST': 	 	context = RequestContext(request) def contacts(request):    	return HttpResponseRedirect('/rango/new1/') 	send_mail(name,query,fromemail,toemail,fail_silently=False)	 	 	toemail=[email] 	fromemail=settings.EMAIL_HOST_USER; 		return render_to_response('contact.html',{'error':error,'name':name,'email':email,'message':query}, context) 		query=request.POST.get('message') 		email=request.POST.get('email') 		name=request.POST.get('name') 	if err == True: 			error.append("please enter message") 			err=True 		if not query: 				error.append("please enter email correctly") 			else: 				error.append("please enter email") 			if not email: 			err=True 		if not email or '@' not in email: 			error.append("please enter name") 			err=True 		if not name:  			query=request.POST.get('message') 		if 'message' in request.POST: 			email=request.POST.get('email') 		if 'email' in request.POST: 			name=request.POST.get('name') 		if 'name' in request.POST: 	if request.method=='POST': 	error=[];	 	err=False 	context = RequestContext(request) 	 def contact1(request):   	return render(request,"contact.html",{}) 	 def contact(request):              return render_to_response('search1.html', context_dict, context) 	context_dict = {'value': sea} 		return render_to_response('search.html', {'error':error}, context) 		error=error[0]	 	if err == True:	 			print error 			error.append('Please enter at most 20 characters.') 			err= True 		elif len(sea)< 3: 			error.append('Enter a search term.') 			err=True 		if not sea: 			sea=request.GET.get('q') 		if 'q' in request.GET: 		 	if request.method=='GET': 	error=[]; 	err=False 	context = RequestContext(request)	 def search1(request):   	return render(request,"search.html",{}) 			 def search(request):            return render(request,"hello.html",context_dict)           context_dict={"var":"god knows wat to do"}  def new1(request):          return render_to_response("hello.html",context_dict,context) 	context_dict={"var":"god knows wat to do"} 	context=RequestContext(request) 	 def new(request):          return JsonResponse({"hi":"how"}) 	 def about1(request):  	return HttpResponse(txt) 	txt="hi rango"+"<a href="+"/rango/>INDEX</a>" def about(request):            	return render_to_response('hello1.html', context_dict, context)         	context_dict = {'page': page_list} 			page_list = Page.objects.filter(category_id=4)		                 else: 			page_list = Page.objects.filter(category_id=3) 		if cat == 'food':         	context = RequestContext(request) 		cat=request.GET.get('category')	         if request.method=='GET': def page(request):  	return render_to_response('hello.html', context_dict, context) 	context_dict = {'categories': category_list} 	print category_list 	category_list = Category.objects.all() 	context = RequestContext(request) def index(request):  # Create your views here.   from django.contrib import auth from rango.forms import * from django.conf import settings from models import * from django.core.mail import send_mail from django.template import RequestContext from django.http import HttpResponse,JsonResponse,HttpResponseRedirect from django.shortcuts import render,render_to_response ad  p  �            �  �  �  J  H  
      �  �  �  �  ~  f  K  0  �  �  �  �  �  O  H  4  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	return render(request, 'loginform.html', {'form': form}) 		form=LoginForm(); 	else: 				return HttpResponseRedirect('/rango/login/') 			else: 				return HttpResponseRedirect('/rango/new1/') 				auth.login(request,user) 			if user is not None: 			user = auth.authenticate(username=Username, password=Password) 			Password=cd['password'] 			Username=cd['username'] 			cd=form.cleaned_data 		if form.is_valid(): 		form=LoginForm(request.POST) 	if request.method=='POST': 	context = RequestContext(request)	 def login(request):  	 	return render(request, 'contactform.html', {'form': form})		 	 		form = ContactForm(initial={'message': 'I love your site!'}) 	else: 			return HttpResponseRedirect('/rango/new1/') 			send_mail(name,message,fromemail,toemail,fail_silently=False) 